--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   13:56:10 10/28/2018
-- Design Name:   
-- Module Name:   C:/Users/Nicolas/Documents/VHDLAtencio/guia04/guiaDeClase04_02_tb.vhd
-- Project Name:  guia04
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: myUartTxTest
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY guiaDeClase04_02_tb IS
END guiaDeClase04_02_tb;
 
ARCHITECTURE behavior OF guiaDeClase04_02_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT myUartTxTest
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         sw : IN  std_logic_vector(3 downto 0);
         tx : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal sw : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal tx : std_logic;

   -- Clock period definitions
   constant clk_period : time := 20 ns;
 
 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: myUartTxTest PORT MAP (
          clk => clk,
          rst => rst,
          sw => sw,
          tx => tx
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin	
		sw<="0000";
		rst<='1';
		wait for 1000 nS;
			
		sw<="1111";
		wait for 100 ns;
		rst<='0';
		wait for clk_period*100000;
		
		sw<="0010";
		wait for clk_period*100000;
		rst<='1';
		wait for 200 ns;
		rst<='0';
		wait;

--		rst<='1';
--		wait for 100 ns;
--		rst<='0';
--		wait for 100 ns;	
--      wait;
   end process;

END;
