--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   15:56:43 10/17/2018
-- Design Name:   
-- Module Name:   C:/Users/Nicolas/Documents/VHDLAtencio/guia02/guiaDeClase02_04_tb.vhd
-- Project Name:  guia02
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: myFFDREN
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY guiaDeClase02_04_tb IS
END guiaDeClase02_04_tb;
 
ARCHITECTURE behavior OF guiaDeClase02_04_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT myFFDREN
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         ena : IN  std_logic;
         d : IN  std_logic_vector(3 downto 0);
         q : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal ena : std_logic := '0';
   signal d : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal q : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant clk_period : time := 100 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: myFFDREN PORT MAP (
          clk => clk,
          rst => rst,
          ena => ena,
          d => d,
          q => q
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
	
		ena<='1';
		rst<='1';
		d<="1111";
		wait for 100 ns;	
		
		ena<='0';
		rst<='0';
		d<="1010";
		wait for 100 ns;	
		d<="1101";
		wait for 100 ns;
      d<="0101";
		wait for 100 ns;	
		d<="1100";
		wait for 100 ns;
      d<="0000";
		wait for 100 ns;	
		d<="0000";
		wait for 100 ns;
      d<="1111";
		wait for 100 ns;	
		d<="1111";
		wait for 100 ns;
		
		
		ena<='0';
		rst<='1';
		d<="1010";
		wait for 100 ns;	
		d<="1101";
		wait for 100 ns;
      d<="0101";
		wait for 100 ns;	
		d<="1100";
		wait for 100 ns;
      d<="0000";
		wait for 100 ns;	
		d<="0000";
		wait for 100 ns;
      d<="1111";
		wait for 100 ns;	
		d<="1111";
		wait for 100 ns;
		
		
		ena<='1';
		rst<='0';
		d<="1010";
		wait for 100 ns;	
		d<="1101";
		wait for 100 ns;
      d<="0101";
		wait for 100 ns;	
		d<="1100";
		wait for 100 ns;
      d<="0000";
		wait for 100 ns;	
		d<="0000";
		wait for 100 ns;
      d<="1111";
		wait for 100 ns;	
		d<="1111";
		wait for 100 ns;
		
		
		ena<='1';
		rst<='1';
		d<="1010";
		wait for 100 ns;	
		d<="1101";
		wait for 100 ns;
      d<="0101";
		wait for 100 ns;	
		d<="1100";
		wait for 100 ns;
      d<="0000";
		wait for 100 ns;	
		d<="0000";
		wait for 100 ns;
      d<="1111";
		wait for 100 ns;	
		d<="1111";
		wait for 100 ns;

		ena<='0';
		rst<='0';
		wait for 100 ns;
	
	
   end process;

END;
