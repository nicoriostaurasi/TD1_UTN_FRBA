----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:37:43 09/28/2018 
-- Design Name: 
-- Module Name:    guiaDeClase00_04 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity guiaDeClase00_04 is
    Port ( a : in  STD_LOGIC_VECTOR (3 downto 0);
           p : out  STD_LOGIC);
end guiaDeClase00_04;

architecture Behavioral of guiaDeClase00_04 is

begin
p<=(a(3) xor a(2)) xor (a(1) xor a(0));
end Behavioral;

